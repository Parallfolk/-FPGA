////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 2013-2021 Efinix Inc. All rights reserved.              
//
// This   document  contains  proprietary information  which   is        
// protected by  copyright. All rights  are reserved.  This notice       
// refers to original work by Efinix, Inc. which may be derivitive       
// of other work distributed under license of the authors.  In the       
// case of derivative work, nothing in this notice overrides the         
// original author's license agreement.  Where applicable, the           
// original license agreement is included in it's original               
// unmodified form immediately below this header.                        
//                                                                       
// WARRANTY DISCLAIMER.                                                  
//     THE  DESIGN, CODE, OR INFORMATION ARE PROVIDED “AS IS” AND        
//     EFINIX MAKES NO WARRANTIES, EXPRESS OR IMPLIED WITH               
//     RESPECT THERETO, AND EXPRESSLY DISCLAIMS ANY IMPLIED WARRANTIES,  
//     INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF          
//     MERCHANTABILITY, NON-INFRINGEMENT AND FITNESS FOR A PARTICULAR    
//     PURPOSE.  SOME STATES DO NOT ALLOW EXCLUSIONS OF AN IMPLIED       
//     WARRANTY, SO THIS DISCLAIMER MAY NOT APPLY TO LICENSEE.           
//                                                                       
// LIMITATION OF LIABILITY.                                              
//     NOTWITHSTANDING ANYTHING TO THE CONTRARY, EXCEPT FOR BODILY       
//     INJURY, EFINIX SHALL NOT BE LIABLE WITH RESPECT TO ANY SUBJECT    
//     MATTER OF THIS AGREEMENT UNDER TORT, CONTRACT, STRICT LIABILITY   
//     OR ANY OTHER LEGAL OR EQUITABLE THEORY (I) FOR ANY INDIRECT,      
//     SPECIAL, INCIDENTAL, EXEMPLARY OR CONSEQUENTIAL DAMAGES OF ANY    
//     CHARACTER INCLUDING, WITHOUT LIMITATION, DAMAGES FOR LOSS OF      
//     GOODWILL, DATA OR PROFIT, WORK STOPPAGE, OR COMPUTER FAILURE OR   
//     MALFUNCTION, OR IN ANY EVENT (II) FOR ANY AMOUNT IN EXCESS, IN    
//     THE AGGREGATE, OF THE FEE PAID BY LICENSEE TO EFINIX HEREUNDER    
//     (OR, IF THE FEE HAS BEEN WAIVED, $100), EVEN IF EFINIX SHALL HAVE 
//     BEEN INFORMED OF THE POSSIBILITY OF SUCH DAMAGES.  SOME STATES DO 
//     NOT ALLOW THE EXCLUSION OR LIMITATION OF INCIDENTAL OR            
//     CONSEQUENTIAL DAMAGES, SO THIS LIMITATION AND EXCLUSION MAY NOT   
//     APPLY TO LICENSEE.                                                
//
////////////////////////////////////////////////////////////////////////////////

    localparam AXI_IF  = 0;
    localparam AXI_DBW = 128;
    localparam AXI_SBW = AXI_DBW/8;
    localparam DDIN_MODE = 0;
    localparam AXI_AWR_DEPTH = 16;
    localparam AXI_R_DEPTH = 256;
    localparam AXI_W_DEPTH = 256;
    localparam CAL_CLK_CH = 4;
    localparam CAL_DQ_STEPS = 8;
    localparam CAL_MODE = 2;
    localparam CAL_RWDS_STEPS = 8;
    localparam CR0_DPD = 1;
    localparam CR0_FLE = 1;
    localparam CR0_ILC = 2;
    localparam CR0_HBE = 1;
    localparam CR0_ODS = 0;
    localparam CR1_HSE = 0;
    localparam CR0_WBL = 3;
    localparam CR1_PAR = 0;
    localparam CR1_MCT = 1;
    localparam RAM_ABW = 25;
    localparam RAM_DBW = 16;
    localparam RDO_DELAY = 3;
    localparam TRH = 200000;
    localparam TRTR = 40000;
    localparam TVCS = 150000000;
    localparam CAL_BYTES = 200;
    localparam MHZ = 200;
    localparam TCSM = 4000000;
	localparam DUAL_RAM = 0;
	localparam INDIVI_DUAL_CAL = 0;
